`timescale 1ns / 1ps

module S_boxes(
	 input rst_n,
    input [0:47] S_in,
    output [0:31] S_out
    );
reg [0:3] s1 [0:3][0:15]; //��ά���飬4��16�У����ݿ��4bit��0~15����
reg [0:3] s2 [0:3][0:15];
reg [0:3] s3 [0:3][0:15];
reg [0:3] s4 [0:3][0:15];
reg [0:3] s5 [0:3][0:15];
reg [0:3] s6 [0:3][0:15];
reg [0:3] s7 [0:3][0:15];
reg [0:3] s8 [0:3][0:15];

wire [0:3] so1,so2,so3,so4,so5,so6,so7,so8;

//s1
always@(negedge rst_n) begin
	s1[0][0]=4'd14; s1[0][1]=4'd4; s1[0][2]=4'd13; s1[0][3]=4'd1; s1[0][4]=4'd2; s1[0][5]=4'd15; s1[0][6]=4'd11; s1[0][7]=4'd8; s1[0][8]=4'd3; s1[0][9]=4'd10; s1[0][10]=4'd6; s1[0][11]=4'd12; s1[0][12]=4'd5; s1[0][13]=4'd9; s1[0][14]=4'd0; s1[0][15]=4'd7; s1[1][0]=4'd0; s1[1][1]=4'd15; s1[1][2]=4'd7; s1[1][3]=4'd4; s1[1][4]=4'd14; s1[1][5]=4'd2; s1[1][6]=4'd13; s1[1][7]=4'd1; s1[1][8]=4'd10; s1[1][9]=4'd6; s1[1][10]=4'd12; s1[1][11]=4'd11; s1[1][12]=4'd9; s1[1][13]=4'd5; s1[1][14]=4'd3; s1[1][15]=4'd8; s1[2][0]=4'd4; s1[2][1]=4'd1; s1[2][2]=4'd14; s1[2][3]=4'd8; s1[2][4]=4'd13; s1[2][5]=4'd6; s1[2][6]=4'd2; s1[2][7]=4'd11; s1[2][8]=4'd15; s1[2][9]=4'd12; s1[2][10]=4'd9; s1[2][11]=4'd7; s1[2][12]=4'd3; s1[2][13]=4'd10; s1[2][14]=4'd5; s1[2][15]=4'd0; s1[3][0]=4'd15; s1[3][1]=4'd12; s1[3][2]=4'd8; s1[3][3]=4'd2; s1[3][4]=4'd4; s1[3][5]=4'd9; s1[3][6]=4'd1; s1[3][7]=4'd7; s1[3][8]=4'd5; s1[3][9]=4'd11; s1[3][10]=4'd3; s1[3][11]=4'd14; s1[3][12]=4'd10; s1[3][13]=4'd0; s1[3][14]=4'd6; s1[3][15]=4'd13;
end

//s2
always@(negedge rst_n) begin
	s2[0][0]=4'd15; s2[0][1]=4'd1; s2[0][2]=4'd8; s2[0][3]=4'd14; s2[0][4]=4'd6; s2[0][5]=4'd11; s2[0][6]=4'd3; s2[0][7]=4'd4; s2[0][8]=4'd9; s2[0][9]=4'd7; s2[0][10]=4'd2; s2[0][11]=4'd13; s2[0][12]=4'd12; s2[0][13]=4'd0; s2[0][14]=4'd5; s2[0][15]=4'd10; s2[1][0]=4'd3; s2[1][1]=4'd13; s2[1][2]=4'd4; s2[1][3]=4'd7; s2[1][4]=4'd15; s2[1][5]=4'd2; s2[1][6]=4'd8; s2[1][7]=4'd14; s2[1][8]=4'd12; s2[1][9]=4'd0; s2[1][10]=4'd1; s2[1][11]=4'd10; s2[1][12]=4'd6; s2[1][13]=4'd9; s2[1][14]=4'd11; s2[1][15]=4'd5; s2[2][0]=4'd0; s2[2][1]=4'd14; s2[2][2]=4'd7; s2[2][3]=4'd11; s2[2][4]=4'd10; s2[2][5]=4'd4; s2[2][6]=4'd13; s2[2][7]=4'd1; s2[2][8]=4'd5; s2[2][9]=4'd8; s2[2][10]=4'd12; s2[2][11]=4'd6; s2[2][12]=4'd9; s2[2][13]=4'd3; s2[2][14]=4'd2; s2[2][15]=4'd15; s2[3][0]=4'd13; s2[3][1]=4'd8; s2[3][2]=4'd10; s2[3][3]=4'd1; s2[3][4]=4'd3; s2[3][5]=4'd15; s2[3][6]=4'd4; s2[3][7]=4'd2; s2[3][8]=4'd11; s2[3][9]=4'd6; s2[3][10]=4'd7; s2[3][11]=4'd12; s2[3][12]=4'd0; s2[3][13]=4'd5; s2[3][14]=4'd14; s2[3][15]=4'd9;
end

//s3
always@(negedge rst_n) begin
	s3[0][0]=4'd10; s3[0][1]=4'd0; s3[0][2]=4'd9; s3[0][3]=4'd14; s3[0][4]=4'd6; s3[0][5]=4'd3; s3[0][6]=4'd15; s3[0][7]=4'd5; s3[0][8]=4'd1; s3[0][9]=4'd13; s3[0][10]=4'd12; s3[0][11]=4'd7; s3[0][12]=4'd11; s3[0][13]=4'd4; s3[0][14]=4'd2; s3[0][15]=4'd8; s3[1][0]=4'd13; s3[1][1]=4'd7; s3[1][2]=4'd0; s3[1][3]=4'd9; s3[1][4]=4'd3; s3[1][5]=4'd4; s3[1][6]=4'd6; s3[1][7]=4'd10; s3[1][8]=4'd2; s3[1][9]=4'd8; s3[1][10]=4'd5; s3[1][11]=4'd14; s3[1][12]=4'd12; s3[1][13]=4'd11; s3[1][14]=4'd15; s3[1][15]=4'd1; s3[2][0]=4'd13; s3[2][1]=4'd6; s3[2][2]=4'd4; s3[2][3]=4'd9; s3[2][4]=4'd8; s3[2][5]=4'd15; s3[2][6]=4'd3; s3[2][7]=4'd0; s3[2][8]=4'd11; s3[2][9]=4'd1; s3[2][10]=4'd2; s3[2][11]=4'd12; s3[2][12]=4'd5; s3[2][13]=4'd10; s3[2][14]=4'd14; s3[2][15]=4'd7; s3[3][0]=4'd1; s3[3][1]=4'd10; s3[3][2]=4'd13; s3[3][3]=4'd0; s3[3][4]=4'd6; s3[3][5]=4'd9; s3[3][6]=4'd8; s3[3][7]=4'd7; s3[3][8]=4'd4; s3[3][9]=4'd15; s3[3][10]=4'd14; s3[3][11]=4'd3; s3[3][12]=4'd11; s3[3][13]=4'd5; s3[3][14]=4'd2; s3[3][15]=4'd12;
end

//s4
always@(negedge rst_n) begin
	s4[0][0]=4'd7; s4[0][1]=4'd13; s4[0][2]=4'd14; s4[0][3]=4'd3; s4[0][4]=4'd0; s4[0][5]=4'd6; s4[0][6]=4'd9; s4[0][7]=4'd10; s4[0][8]=4'd1; s4[0][9]=4'd2; s4[0][10]=4'd8; s4[0][11]=4'd5; s4[0][12]=4'd11; s4[0][13]=4'd12; s4[0][14]=4'd4; s4[0][15]=4'd15; s4[1][0]=4'd13; s4[1][1]=4'd8; s4[1][2]=4'd11; s4[1][3]=4'd5; s4[1][4]=4'd6; s4[1][5]=4'd15; s4[1][6]=4'd0; s4[1][7]=4'd3; s4[1][8]=4'd4; s4[1][9]=4'd7; s4[1][10]=4'd2; s4[1][11]=4'd12; s4[1][12]=4'd1; s4[1][13]=4'd10; s4[1][14]=4'd14; s4[1][15]=4'd9; s4[2][0]=4'd10; s4[2][1]=4'd6; s4[2][2]=4'd9; s4[2][3]=4'd0; s4[2][4]=4'd12; s4[2][5]=4'd11; s4[2][6]=4'd7; s4[2][7]=4'd13; s4[2][8]=4'd15; s4[2][9]=4'd1; s4[2][10]=4'd3; s4[2][11]=4'd14; s4[2][12]=4'd5; s4[2][13]=4'd2; s4[2][14]=4'd8; s4[2][15]=4'd4; s4[3][0]=4'd3; s4[3][1]=4'd15; s4[3][2]=4'd0; s4[3][3]=4'd6; s4[3][4]=4'd10; s4[3][5]=4'd1; s4[3][6]=4'd13; s4[3][7]=4'd8; s4[3][8]=4'd9; s4[3][9]=4'd4; s4[3][10]=4'd5; s4[3][11]=4'd11; s4[3][12]=4'd12; s4[3][13]=4'd7; s4[3][14]=4'd2; s4[3][15]=4'd14;
end

//s5
always@(negedge rst_n) begin
	s5[0][0]=4'd2; s5[0][1]=4'd12; s5[0][2]=4'd4; s5[0][3]=4'd1; s5[0][4]=4'd7; s5[0][5]=4'd10; s5[0][6]=4'd11; s5[0][7]=4'd6; s5[0][8]=4'd8; s5[0][9]=4'd5; s5[0][10]=4'd3; s5[0][11]=4'd15; s5[0][12]=4'd13; s5[0][13]=4'd0; s5[0][14]=4'd14; s5[0][15]=4'd9; s5[1][0]=4'd14; s5[1][1]=4'd11; s5[1][2]=4'd2; s5[1][3]=4'd12; s5[1][4]=4'd4; s5[1][5]=4'd7; s5[1][6]=4'd13; s5[1][7]=4'd1; s5[1][8]=4'd5; s5[1][9]=4'd0; s5[1][10]=4'd15; s5[1][11]=4'd10; s5[1][12]=4'd3; s5[1][13]=4'd9; s5[1][14]=4'd8; s5[1][15]=4'd6; s5[2][0]=4'd4; s5[2][1]=4'd2; s5[2][2]=4'd1; s5[2][3]=4'd11; s5[2][4]=4'd10; s5[2][5]=4'd13; s5[2][6]=4'd7; s5[2][7]=4'd8; s5[2][8]=4'd15; s5[2][9]=4'd9; s5[2][10]=4'd12; s5[2][11]=4'd5; s5[2][12]=4'd6; s5[2][13]=4'd3; s5[2][14]=4'd0; s5[2][15]=4'd14; s5[3][0]=4'd11; s5[3][1]=4'd8; s5[3][2]=4'd12; s5[3][3]=4'd7; s5[3][4]=4'd1; s5[3][5]=4'd14; s5[3][6]=4'd2; s5[3][7]=4'd13; s5[3][8]=4'd6; s5[3][9]=4'd15; s5[3][10]=4'd0; s5[3][11]=4'd9; s5[3][12]=4'd10; s5[3][13]=4'd4; s5[3][14]=4'd5; s5[3][15]=4'd3;
end

//s6
always@(negedge rst_n) begin
	s6[0][0]=4'd12; s6[0][1]=4'd1; s6[0][2]=4'd10; s6[0][3]=4'd15; s6[0][4]=4'd9; s6[0][5]=4'd2; s6[0][6]=4'd6; s6[0][7]=4'd8; s6[0][8]=4'd0; s6[0][9]=4'd13; s6[0][10]=4'd3; s6[0][11]=4'd4; s6[0][12]=4'd14; s6[0][13]=4'd7; s6[0][14]=4'd5; s6[0][15]=4'd11; s6[1][0]=4'd10; s6[1][1]=4'd15; s6[1][2]=4'd4; s6[1][3]=4'd2; s6[1][4]=4'd7; s6[1][5]=4'd12; s6[1][6]=4'd9; s6[1][7]=4'd5; s6[1][8]=4'd6; s6[1][9]=4'd1; s6[1][10]=4'd13; s6[1][11]=4'd14; s6[1][12]=4'd0; s6[1][13]=4'd11; s6[1][14]=4'd3; s6[1][15]=4'd8; s6[2][0]=4'd9; s6[2][1]=4'd14; s6[2][2]=4'd15; s6[2][3]=4'd5; s6[2][4]=4'd2; s6[2][5]=4'd8; s6[2][6]=4'd12; s6[2][7]=4'd3; s6[2][8]=4'd7; s6[2][9]=4'd0; s6[2][10]=4'd4; s6[2][11]=4'd10; s6[2][12]=4'd1; s6[2][13]=4'd13; s6[2][14]=4'd11; s6[2][15]=4'd6; s6[3][0]=4'd4; s6[3][1]=4'd3; s6[3][2]=4'd2; s6[3][3]=4'd12; s6[3][4]=4'd9; s6[3][5]=4'd5; s6[3][6]=4'd15; s6[3][7]=4'd10; s6[3][8]=4'd11; s6[3][9]=4'd14; s6[3][10]=4'd1; s6[3][11]=4'd7; s6[3][12]=4'd6; s6[3][13]=4'd0; s6[3][14]=4'd8; s6[3][15]=4'd13;
end

//s7
always@(negedge rst_n) begin
	s7[0][0]=4'd4; s7[0][1]=4'd11; s7[0][2]=4'd2; s7[0][3]=4'd14; s7[0][4]=4'd15; s7[0][5]=4'd0; s7[0][6]=4'd8; s7[0][7]=4'd13; s7[0][8]=4'd3; s7[0][9]=4'd12; s7[0][10]=4'd9; s7[0][11]=4'd7; s7[0][12]=4'd5; s7[0][13]=4'd10; s7[0][14]=4'd6; s7[0][15]=4'd1; s7[1][0]=4'd13; s7[1][1]=4'd0; s7[1][2]=4'd11; s7[1][3]=4'd7; s7[1][4]=4'd4; s7[1][5]=4'd9; s7[1][6]=4'd1; s7[1][7]=4'd10; s7[1][8]=4'd14; s7[1][9]=4'd3; s7[1][10]=4'd5; s7[1][11]=4'd12; s7[1][12]=4'd2; s7[1][13]=4'd15; s7[1][14]=4'd8; s7[1][15]=4'd6; s7[2][0]=4'd1; s7[2][1]=4'd4; s7[2][2]=4'd11; s7[2][3]=4'd13; s7[2][4]=4'd12; s7[2][5]=4'd3; s7[2][6]=4'd7; s7[2][7]=4'd14; s7[2][8]=4'd10; s7[2][9]=4'd15; s7[2][10]=4'd6; s7[2][11]=4'd8; s7[2][12]=4'd0; s7[2][13]=4'd5; s7[2][14]=4'd9; s7[2][15]=4'd2; s7[3][0]=4'd6; s7[3][1]=4'd11; s7[3][2]=4'd13; s7[3][3]=4'd8; s7[3][4]=4'd1; s7[3][5]=4'd4; s7[3][6]=4'd10; s7[3][7]=4'd7; s7[3][8]=4'd9; s7[3][9]=4'd5; s7[3][10]=4'd0; s7[3][11]=4'd15; s7[3][12]=4'd14; s7[3][13]=4'd2; s7[3][14]=4'd3; s7[3][15]=4'd12;
end

//s8
always@(negedge rst_n) begin
	s8[0][0]=4'd13; s8[0][1]=4'd2; s8[0][2]=4'd8; s8[0][3]=4'd4; s8[0][4]=4'd6; s8[0][5]=4'd15; s8[0][6]=4'd11; s8[0][7]=4'd1; s8[0][8]=4'd10; s8[0][9]=4'd9; s8[0][10]=4'd3; s8[0][11]=4'd14; s8[0][12]=4'd5; s8[0][13]=4'd0; s8[0][14]=4'd12; s8[0][15]=4'd7; s8[1][0]=4'd1; s8[1][1]=4'd15; s8[1][2]=4'd13; s8[1][3]=4'd8; s8[1][4]=4'd10; s8[1][5]=4'd3; s8[1][6]=4'd7; s8[1][7]=4'd4; s8[1][8]=4'd12; s8[1][9]=4'd5; s8[1][10]=4'd6; s8[1][11]=4'd11; s8[1][12]=4'd0; s8[1][13]=4'd14; s8[1][14]=4'd9; s8[1][15]=4'd2; s8[2][0]=4'd7; s8[2][1]=4'd11; s8[2][2]=4'd4; s8[2][3]=4'd1; s8[2][4]=4'd9; s8[2][5]=4'd12; s8[2][6]=4'd14; s8[2][7]=4'd2; s8[2][8]=4'd0; s8[2][9]=4'd6; s8[2][10]=4'd10; s8[2][11]=4'd13; s8[2][12]=4'd15; s8[2][13]=4'd3; s8[2][14]=4'd5; s8[2][15]=4'd8; s8[3][0]=4'd2; s8[3][1]=4'd1; s8[3][2]=4'd14; s8[3][3]=4'd7; s8[3][4]=4'd4; s8[3][5]=4'd10; s8[3][6]=4'd8; s8[3][7]=4'd13; s8[3][8]=4'd15; s8[3][9]=4'd12; s8[3][10]=4'd9; s8[3][11]=4'd0; s8[3][12]=4'd3; s8[3][13]=4'd5; s8[3][14]=4'd6; s8[3][15]=4'd11;
end

assign so1 = s1[{S_in[0],S_in[5]}][S_in[1:4]];
assign so2 = s2[{S_in[6],S_in[11]}][S_in[7:10]];
assign so3 = s3[{S_in[12],S_in[17]}][S_in[13:16]];
assign so4 = s4[{S_in[18],S_in[23]}][S_in[19:22]];
assign so5 = s5[{S_in[24],S_in[29]}][S_in[25:28]];
assign so6 = s6[{S_in[30],S_in[35]}][S_in[31:34]];
assign so7 = s7[{S_in[36],S_in[41]}][S_in[37:40]];
assign so8 = s8[{S_in[42],S_in[47]}][S_in[43:46]];

assign S_out = {so1,so2,so3,so4,so5,so6,so7,so8};
endmodule


